module self_fifo

end